module ProjectB();


endmodule
